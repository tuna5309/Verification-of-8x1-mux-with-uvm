interface mux_intf();
logic d0;
logic d1;
logic d2;
logic d3;
logic d4;
logic d5;
logic d6;
logic d7;
logic  [2:0] sel; 
logic  out;
endinterface
